magic
tech sky130A
magscale 1 2
timestamp 1725617993
<< locali >>
rect 19047 5685 19253 5691
rect 17586 5652 17770 5658
rect 16107 5595 16305 5601
rect 16107 5409 16113 5595
rect 16299 5409 16305 5595
rect 16107 2397 16305 5409
rect 17586 5480 17592 5652
rect 17764 5480 17770 5652
rect 17586 2434 17770 5480
rect 19047 5491 19053 5685
rect 19247 5491 19253 5685
rect 19047 2661 19253 5491
<< viali >>
rect 16113 5409 16299 5595
rect 16107 2199 16305 2397
rect 17592 5480 17764 5652
rect 19053 5491 19247 5685
rect 19047 2455 19253 2661
rect 17586 2250 17770 2434
<< metal1 >>
rect 14102 27654 14108 27846
rect 14300 27654 20724 27846
rect 16104 23796 20724 24000
rect 16104 13384 16308 23796
rect 27266 22454 27466 25036
rect 17586 21852 20756 22036
rect 16107 5595 16305 13384
rect 17586 5658 17770 21852
rect 19047 20242 20853 20448
rect 19047 5685 19253 20242
rect 16107 5409 16113 5595
rect 16299 5409 16305 5595
rect 17580 5652 17776 5658
rect 17580 5480 17592 5652
rect 17764 5480 17776 5652
rect 17580 5474 17776 5480
rect 19047 5491 19053 5685
rect 19247 5491 19253 5685
rect 19047 5479 19253 5491
rect 16107 5397 16305 5409
rect 15127 3237 15356 3243
rect 15356 3008 20888 3237
rect 15127 3002 15356 3008
rect 19035 2661 19265 2667
rect 19035 2455 19047 2661
rect 19253 2584 26675 2661
rect 27268 2634 27464 22454
rect 19253 2455 26678 2584
rect 19035 2449 19265 2455
rect 17574 2434 17782 2440
rect 16095 2397 16317 2403
rect 16095 2199 16107 2397
rect 16305 2199 16317 2397
rect 17574 2250 17586 2434
rect 17770 2250 17782 2434
rect 17574 2244 17782 2250
rect 16095 2193 16317 2199
rect 16107 1359 16305 2193
rect 17586 2066 17770 2244
rect 17586 2020 22790 2066
rect 17586 1882 22814 2020
rect 16107 1350 18814 1359
rect 16107 1162 18950 1350
rect 16107 1161 16305 1162
rect 18770 852 18950 1162
rect 22634 1026 22814 1882
rect 26498 1176 26678 2455
rect 27268 2438 30544 2634
rect 30362 1306 30542 2438
rect 18764 672 18770 852
rect 18950 672 18956 852
rect 22628 846 22634 1026
rect 22814 846 22820 1026
rect 26492 996 26498 1176
rect 26678 996 26684 1176
rect 30356 1126 30362 1306
rect 30542 1126 30548 1306
<< via1 >>
rect 14108 27654 14300 27846
rect 15127 3008 15356 3237
rect 18770 672 18950 852
rect 22634 846 22814 1026
rect 26498 996 26678 1176
rect 30362 1126 30542 1306
<< metal2 >>
rect 14108 27846 14300 27852
rect 13673 27654 13682 27846
rect 13874 27654 14108 27846
rect 14108 27648 14300 27654
rect 14380 3237 14599 3241
rect 14375 3232 15127 3237
rect 14375 3013 14380 3232
rect 14599 3013 15127 3232
rect 14375 3008 15127 3013
rect 15356 3008 15362 3237
rect 14380 3004 14599 3008
rect 30362 1306 30542 1312
rect 26498 1176 26678 1182
rect 22634 1026 22814 1032
rect 18770 852 18950 858
rect 30362 1021 30542 1126
rect 26498 891 26678 996
rect 22634 825 22814 846
rect 18770 653 18950 672
rect 22630 655 22639 825
rect 22809 655 22818 825
rect 26494 721 26503 891
rect 26673 721 26682 891
rect 30358 851 30367 1021
rect 30537 851 30546 1021
rect 30362 846 30542 851
rect 26498 716 26678 721
rect 18766 483 18775 653
rect 18945 483 18954 653
rect 22634 650 22814 655
rect 18770 478 18950 483
<< via2 >>
rect 13682 27654 13874 27846
rect 14380 3013 14599 3232
rect 22639 655 22809 825
rect 26503 721 26673 891
rect 30367 851 30537 1021
rect 18775 483 18945 653
<< metal3 >>
rect 13677 27846 13879 27851
rect 13208 27654 13214 27846
rect 13406 27654 13682 27846
rect 13874 27654 13879 27846
rect 13677 27649 13879 27654
rect 13784 3237 14011 3242
rect 13783 3236 14604 3237
rect 13783 3009 13784 3236
rect 14011 3232 14604 3236
rect 14011 3013 14380 3232
rect 14599 3013 14604 3232
rect 14011 3009 14604 3013
rect 13783 3008 14604 3009
rect 13784 3003 14011 3008
rect 30362 1021 30542 1026
rect 26498 891 26678 896
rect 22634 825 22814 830
rect 18770 653 18950 658
rect 18770 483 18775 653
rect 18945 483 18950 653
rect 18770 419 18950 483
rect 22634 655 22639 825
rect 22809 655 22814 825
rect 22634 591 22814 655
rect 26498 721 26503 891
rect 26673 721 26678 891
rect 26498 613 26678 721
rect 30362 851 30367 1021
rect 30537 851 30542 1021
rect 30362 679 30542 851
rect 18765 241 18771 419
rect 18949 241 18955 419
rect 22634 413 22635 591
rect 22813 413 22814 591
rect 26493 435 26499 613
rect 26677 435 26683 613
rect 30357 501 30363 679
rect 30541 501 30547 679
rect 30362 500 30542 501
rect 26498 434 26678 435
rect 22634 412 22814 413
rect 22635 407 22813 412
rect 18770 240 18950 241
<< via3 >>
rect 13214 27654 13406 27846
rect 13784 3009 14011 3236
rect 18771 241 18949 419
rect 22635 413 22813 591
rect 26499 435 26677 613
rect 30363 501 30541 679
<< metal4 >>
rect 6134 44190 6194 45152
rect 6686 44190 6746 45152
rect 7238 44190 7298 45152
rect 7790 44190 7850 45152
rect 8342 44190 8402 45152
rect 8894 44190 8954 45152
rect 9446 44190 9506 45152
rect 9998 44190 10058 45152
rect 10550 44190 10610 45152
rect 11102 44190 11162 45152
rect 11654 44190 11714 45152
rect 12206 44190 12266 45152
rect 12758 44190 12818 45152
rect 13310 44190 13370 45152
rect 13862 44190 13922 45152
rect 14414 44190 14474 45152
rect 14966 44190 15026 45152
rect 15518 44190 15578 45152
rect 16070 44190 16130 45152
rect 16622 44190 16682 45152
rect 17174 44190 17234 45152
rect 17726 44190 17786 45152
rect 18278 44190 18338 45152
rect 18830 44190 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 803 44152 18994 44190
rect 200 27943 600 44152
rect 800 43800 18994 44152
rect 200 27558 244 27943
rect 200 1000 600 27558
rect 800 22776 1200 43800
rect 18604 43762 18994 43800
rect 3498 27534 3518 27967
rect 3961 27846 12889 27967
rect 13213 27846 13407 27847
rect 3961 27654 13214 27846
rect 13406 27654 13407 27846
rect 3961 27534 12889 27654
rect 13213 27653 13407 27654
rect 800 22376 3510 22776
rect 800 3322 1200 22376
rect 800 3237 13452 3322
rect 800 3236 14012 3237
rect 800 3009 13784 3236
rect 14011 3009 14012 3236
rect 800 3008 14012 3009
rect 800 2922 13452 3008
rect 800 1000 1200 2922
rect 30362 679 30542 680
rect 26498 613 26678 614
rect 22634 591 22814 592
rect 18770 419 18950 420
rect 18770 241 18771 419
rect 18949 241 18950 419
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 241
rect 22634 413 22635 591
rect 22813 413 22814 591
rect 22634 0 22814 413
rect 26498 435 26499 613
rect 26677 435 26678 613
rect 26498 0 26678 435
rect 30362 501 30363 679
rect 30541 501 30542 679
rect 30362 0 30542 501
<< via4 >>
rect 244 27558 629 27943
rect 3518 27534 3961 27967
<< metal5 >>
rect 3494 27967 3985 27991
rect 220 27943 3518 27967
rect 220 27558 244 27943
rect 629 27558 3518 27943
rect 220 27534 3518 27558
rect 3961 27534 3985 27967
rect 3494 27510 3985 27534
use ota5t_1  ota5t_1_0
timestamp 1723807770
transform 1 0 20588 0 1 25366
box -24 -22352 6878 2494
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
