magic
tech sky130A
magscale 1 2
timestamp 1723805434
<< viali >>
rect 1276 1112 1462 1146
rect 2740 1112 2932 1146
rect 1166 -2536 1316 -2496
rect 2650 -2560 2800 -2508
rect 1250 -5718 1608 -5672
rect 2694 -5684 3042 -5646
<< metal1 >>
rect -6 2294 6726 2494
rect 1180 1146 1549 2294
rect 1180 1112 1276 1146
rect 1462 1112 1549 1146
rect 1180 1104 1549 1112
rect 946 509 1212 944
rect 738 243 1212 509
rect 741 -410 848 243
rect 946 64 1212 243
rect 1580 640 1852 868
rect 2018 640 2182 2294
rect 2645 1146 3008 2294
rect 2645 1112 2740 1146
rect 2932 1112 3008 1146
rect 2645 1099 3008 1112
rect 1580 434 2182 640
rect 1580 342 1848 434
rect 1580 152 1852 342
rect 2414 328 2668 944
rect 2232 196 2668 328
rect 1339 -410 1501 -63
rect 741 -572 1847 -410
rect 2009 -572 2015 -410
rect -24 -1556 256 -1356
rect 456 -1556 462 -1356
rect 741 -2102 848 -572
rect 2232 -858 2364 196
rect 2414 64 2668 196
rect 3046 643 3312 950
rect 3494 643 3673 2294
rect 6078 1952 6576 2046
rect 6072 1848 6078 1952
rect 6182 1942 6576 1952
rect 6182 1848 6188 1942
rect 3046 421 3673 643
rect 3046 377 3579 421
rect 3046 90 3312 377
rect 2714 -398 2888 -79
rect 6472 -366 6576 1942
rect 2415 -410 2577 -404
rect 2714 -410 2900 -398
rect 2577 -560 2900 -410
rect 6472 -558 6878 -366
rect 2577 -572 2889 -560
rect 2415 -578 2577 -572
rect 6472 -858 6576 -558
rect 6678 -852 6878 -558
rect 2232 -990 6576 -858
rect 2232 -1200 2364 -990
rect 2232 -1338 2364 -1332
rect 938 -1356 1138 -1350
rect 1138 -1554 1286 -1356
rect 938 -1562 1188 -1554
rect 1232 -1585 1286 -1554
rect 1232 -1656 1289 -1585
rect 1239 -1925 1289 -1656
rect 1668 -1724 3516 -1536
rect 1304 -2084 1492 -1964
rect 1668 -2084 1856 -1724
rect 741 -2209 1195 -2102
rect 1304 -2272 1856 -2084
rect 2482 -2136 2668 -1988
rect 2226 -2268 2232 -2136
rect 2364 -2268 2668 -2136
rect 1304 -2346 1492 -2272
rect 1686 -2483 1839 -2272
rect 2482 -2380 2668 -2268
rect 2780 -2058 2982 -1988
rect 3328 -2058 3516 -1724
rect 2780 -2246 3516 -2058
rect 2780 -2376 2982 -2246
rect 3655 -2409 3661 -2361
rect 2667 -2443 3661 -2409
rect 1139 -2496 1349 -2485
rect 1139 -2536 1166 -2496
rect 1316 -2536 1349 -2496
rect 1139 -2842 1349 -2536
rect 3655 -2492 3661 -2443
rect 3792 -2492 3798 -2361
rect 1686 -2642 1839 -2636
rect 2620 -2508 2830 -2493
rect 2620 -2560 2650 -2508
rect 2800 -2560 2830 -2508
rect 2620 -2842 2830 -2560
rect 1139 -3052 3583 -2842
rect 0 -3528 2968 -3328
rect 3168 -3528 3174 -3328
rect 1680 -3852 1686 -3699
rect 1839 -3852 2041 -3699
rect 2194 -3852 2200 -3699
rect 752 -4418 2864 -4362
rect 6 -4927 206 -4916
rect 752 -4927 808 -4418
rect 1406 -4506 1462 -4418
rect 1402 -4554 1462 -4506
rect 1402 -4650 1458 -4554
rect 1236 -4706 1640 -4650
rect 2808 -4672 2864 -4418
rect 6 -5008 808 -4927
rect 3373 -4971 3583 -3052
rect 6 -5064 1214 -5008
rect 6 -5105 807 -5064
rect 6 -5116 206 -5105
rect 2063 -5146 2069 -5050
rect 2165 -5146 2658 -5050
rect 3045 -5181 3583 -4971
rect 1650 -5538 2110 -5338
rect 1214 -5672 1662 -5666
rect 1214 -5718 1250 -5672
rect 1608 -5718 1662 -5672
rect 1214 -5860 1662 -5718
rect 1284 -6174 1484 -5860
rect 1910 -6174 2110 -5538
rect 2644 -5646 3102 -5640
rect 2644 -5684 2694 -5646
rect 3042 -5684 3102 -5646
rect 2644 -5868 3102 -5684
rect 1284 -6374 2110 -6174
rect 1284 -22152 1484 -6374
rect 2772 -22152 2972 -5868
rect 3373 -22152 3583 -5181
rect 5264 -21698 5368 -21692
rect 5368 -21802 5516 -21698
rect 5264 -21808 5368 -21802
rect 5412 -22152 5516 -21802
rect -10 -22352 6442 -22152
<< via1 >>
rect 1847 -572 2009 -410
rect 256 -1556 456 -1356
rect 6078 1848 6182 1952
rect 2415 -572 2577 -410
rect 2232 -1332 2364 -1200
rect 938 -1554 1138 -1356
rect 2232 -2268 2364 -2136
rect 1686 -2636 1839 -2483
rect 3661 -2492 3792 -2361
rect 2968 -3528 3168 -3328
rect 1686 -3852 1839 -3699
rect 2041 -3852 2194 -3699
rect 2069 -5146 2165 -5050
rect 5264 -21802 5368 -21698
<< metal2 >>
rect 6078 1952 6182 1958
rect 6074 1848 6078 1857
rect 6182 1848 6186 1857
rect 6074 1763 6083 1848
rect 6177 1763 6186 1848
rect 6078 1758 6182 1763
rect 1847 -410 2009 -404
rect 2009 -572 2415 -410
rect 2577 -572 2583 -410
rect 1847 -578 2009 -572
rect 2226 -1332 2232 -1200
rect 2364 -1332 2370 -1200
rect 256 -1356 456 -1350
rect 456 -1554 938 -1356
rect 1138 -1554 1144 -1356
rect 456 -1556 880 -1554
rect 256 -1562 456 -1556
rect 2232 -2136 2364 -1332
rect 2232 -2274 2364 -2268
rect 3661 -2361 3792 -2355
rect 1680 -2636 1686 -2483
rect 1839 -2636 1845 -2483
rect 1686 -3699 1839 -2636
rect 2968 -3328 3168 -3322
rect 3661 -3328 3792 -2492
rect 3168 -3528 3792 -3328
rect 2968 -3534 3168 -3528
rect 1686 -3858 1839 -3852
rect 2041 -3699 2194 -3693
rect 2041 -3858 2194 -3852
rect 2069 -5050 2165 -3858
rect 2069 -5152 2165 -5146
rect 5119 -21698 5213 -21694
rect 5114 -21703 5264 -21698
rect 5114 -21797 5119 -21703
rect 5213 -21797 5264 -21703
rect 5114 -21802 5264 -21797
rect 5368 -21802 5374 -21698
rect 5119 -21806 5213 -21802
<< via2 >>
rect 6083 1848 6177 1857
rect 6083 1763 6177 1848
rect 5119 -21797 5213 -21703
<< metal3 >>
rect 6078 1857 6182 1862
rect 6078 1763 6083 1857
rect 6177 1763 6182 1857
rect 6078 1743 6182 1763
rect 6078 1641 6079 1743
rect 6181 1641 6182 1743
rect 6078 1640 6182 1641
rect 6079 1635 6181 1640
rect 4978 -21699 5218 -21698
rect 4973 -21801 4979 -21699
rect 5081 -21703 5218 -21699
rect 5081 -21797 5119 -21703
rect 5213 -21797 5218 -21703
rect 5081 -21801 5218 -21797
rect 4978 -21802 5218 -21801
<< via3 >>
rect 6079 1641 6181 1743
rect 4979 -21801 5081 -21699
<< metal4 >>
rect 6078 1743 6362 1744
rect 6078 1641 6079 1743
rect 6181 1641 6362 1743
rect 6078 1640 6362 1641
rect 6258 1422 6362 1640
rect 4978 -21699 5082 -21570
rect 4978 -21801 4979 -21699
rect 5081 -21801 5082 -21699
rect 4978 -21802 5082 -21801
use sky130_fd_pr__cap_mim_m3_1_72JAQ7  XC1
timestamp 1723797800
transform 1 0 5176 0 1 -10074
box -1186 -11600 1186 11600
use sky130_fd_pr__nfet_01v8_AHRV9L  XM1
timestamp 1723797800
transform 1 0 2848 0 1 -5100
box -396 -610 396 610
use sky130_fd_pr__pfet_01v8_lvt_GWNSVV  XM2
timestamp 1723797800
transform 1 0 1418 0 1 463
box -396 -719 396 719
use sky130_fd_pr__nfet_01v8_AHRV9L  XM3
timestamp 1723797800
transform 1 0 1434 0 1 -5134
box -396 -610 396 610
use sky130_fd_pr__nfet_01v8_lvt_8TEWK3  XM4
timestamp 1723797800
transform 1 0 2730 0 1 -2174
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_lvt_8TEWK3  XM6
timestamp 1723797800
transform 1 0 1250 0 1 -2158
box -246 -410 246 410
use sky130_fd_pr__pfet_01v8_lvt_GWNSVV  XM7
timestamp 1723797800
transform 1 0 2864 0 1 463
box -396 -719 396 719
<< labels >>
flabel metal1 -6 2294 194 2494 0 FreeSans 256 0 0 0 VCC
port 0 nsew
flabel metal1 -10 -22352 190 -22152 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 0 -3528 200 -3328 0 FreeSans 256 0 0 0 MINUS
port 3 nsew
flabel metal1 6 -5116 206 -4916 0 FreeSans 256 0 0 0 BIAS
port 2 nsew
flabel metal1 -24 -1556 176 -1356 0 FreeSans 256 0 0 0 PLUS
port 4 nsew
flabel metal1 6678 -852 6878 -652 0 FreeSans 256 0 0 0 DIFFOUT
port 1 nsew
flabel metal1 741 -572 1847 -410 0 FreeSans 1600 0 0 0 Vleft
<< end >>
